module led7seg (ILED,SA);
    input [3:0]a;
    output [7:0]LED,SA;

    assign  SA = 4'bZZZ0;
    assign  LED[0] = ;
    assign  LED[1] = ;
    assign  LED[2] = ;
    assign  LED[3] = ;
    assign  LED[4] = ;
    assign  LED[5] = ;
    assign  LED[6] = ;
    assign  LED[7] = 1'b1;
endmodule
