module my_xor ( A, B, Y);
    input A, B;
    output Y;
    
    assign Y = A ^ B;
endmodule